`timescale 1ns / 1ps

module ProcessKey(output reg [48:1] k1,k2,k3,k4,k5,k6,k7,k8,k9,k10,k11,k12,k13,k14,k15,k16,input [64:1] key);
  
  function [56:1] PC1_perm(input [64:1] key);
    integer PC1[56:1];
    integer i;
    reg [56:1] temp_perm;
    begin
			PC1[1] = 57;PC1[2] = 49;PC1[3] = 41;PC1[4] = 33;PC1[5] = 25;PC1[6] = 17;PC1[7] = 9;PC1[8] = 1;PC1[9] = 58;PC1[10] = 50;PC1[11] = 42;PC1[12] = 34;PC1[13] = 26;PC1[14] = 18;PC1[15] = 10;PC1[16] = 2;PC1[17] = 59;PC1[18] = 51;PC1[19] = 43;PC1[20] = 35;PC1[21] = 27;PC1[22] = 19;PC1[23] = 11;PC1[24] = 3;PC1[25] = 60;PC1[26] = 52;PC1[27] = 44;PC1[28] = 36;PC1[29] = 63;PC1[30] = 55;PC1[31] = 47;PC1[32] = 39;PC1[33] = 31;PC1[34] = 23;PC1[35] = 15;PC1[36] = 7;PC1[37] = 62;PC1[38] = 54;PC1[39] = 46;PC1[40] = 38;PC1[41] = 30;PC1[42] = 22;PC1[43] = 14;PC1[44] = 6;PC1[45] = 61;PC1[46] = 53;PC1[47] = 45;PC1[48] = 37;PC1[49] = 29;PC1[50] = 21;PC1[51] = 13;PC1[52] = 5;PC1[53] = 28;PC1[54] = 20;PC1[55] = 12;PC1[56] = 4;
			
			for(i=1; i<=56; i=i+1)
        temp_perm[56-i+1] = key[64-PC1[i]+1];
			
			PC1_perm = temp_perm;
    end
  endfunction
  
  function [48:1] PC2_perm(input [56:1] key_s);
    integer PC2[48:1];
    integer i;
    reg [48:1] temp_perm;
    begin
		PC2[1] = 14;PC2[2] = 17;PC2[3] = 11;PC2[4] = 24;PC2[5] = 1;PC2[6] = 5;PC2[7] = 3;PC2[8] = 28;PC2[9] = 15;PC2[10] = 6;PC2[11] = 21;PC2[12] = 10;PC2[13] = 23;PC2[14] = 19;PC2[15] = 12;PC2[16] = 4;PC2[17] = 26;PC2[18] = 8;PC2[19] = 16;PC2[20] = 7;PC2[21] = 27;PC2[22] = 20;PC2[23] = 13;PC2[24] = 2;PC2[25] = 41;PC2[26] = 52;PC2[27] = 31;PC2[28] = 37;PC2[29] = 47;PC2[30] = 55;PC2[31] = 30;PC2[32] = 40;PC2[33] = 51;PC2[34] = 45;PC2[35] = 33;PC2[36] = 48;PC2[37] = 44;PC2[38] = 49;PC2[39] = 39;PC2[40] = 56;PC2[41] = 34;PC2[42] = 53;PC2[43] = 46;PC2[44] = 42;PC2[45] = 50;PC2[46] = 36;PC2[47] = 29;PC2[48] = 32;
			
			for(i=1; i<=48; i=i+1)
        temp_perm[48-i+1] = key_s[56-PC2[i]+1];

			PC2_perm = temp_perm;
    end
  endfunction

  function [56:1] C_i_D_i(input integer i, input [28:1] C_last, D_last);
    integer shift_left[1:16];
    begin
      shift_left[1] = 1;
      shift_left[2] = 1;
      shift_left[3] = 2;
      shift_left[4] = 2;
      shift_left[5] = 2;
      shift_left[6] = 2;
      shift_left[7] = 2;
      shift_left[8] = 2;
      shift_left[9] = 1;
      shift_left[10] = 2;
      shift_left[11] = 2;
      shift_left[12] = 2;
      shift_left[13] = 2;
      shift_left[14] = 2;
      shift_left[15] = 2;
      shift_left[16] = 1;
      
      if(shift_left[i] == 'd1)
        C_i_D_i = {C_last[27:1], C_last[28], D_last[27:1], D_last[28]};
      else if(shift_left[i] == 'd2)
        C_i_D_i = {C_last[26:1], C_last[28:27], D_last[26:1], D_last[28:27]};
      
    end
  endfunction

  reg [56:1] temp_pc1;
  reg [28:1] C[16:0], D[16:0];
  reg [48:1] K[1:16];
  integer i;
  
  always @(key)
  begin
    temp_pc1 = PC1_perm(key);
    C[0] = temp_pc1[56:29];
    D[0] = temp_pc1[28:1];
    for(i=1; i<=16; i=i+1)
    begin
      {C[i], D[i]} = C_i_D_i(i, C[i-1], D[i-1]);
      K[i] = PC2_perm({C[i], D[i]});
    end
    
    k1 = K[1];
    k2 = K[2];
    k3 = K[3];
    k4 = K[4];
    k5 = K[5];
    k6 = K[6];
    k7 = K[7];
    k8 = K[8];
    k9 = K[9];
    k10 = K[10];
    k11 = K[11];
    k12 = K[12];
    k13 = K[13];
    k14 = K[14];
    k15 = K[15];
    k16 = K[16];
  end
endmodule

module enigma(img,key,enigma);
       input [64:1] img;
       input [64:1] key;
       output reg [64:1] enigma;
       

       function [64:1] IPerm(input [64:1] img);
        integer IP[64:1];
        reg [64:1] z;
        integer i;
              begin
                     IP[1] = 40;
			IP[2] = 8;
			IP[3] = 48;
			IP[4] = 16;
			IP[5] = 56;
			IP[6] = 24;
			IP[7] = 64;
			IP[8] = 32;
			IP[9] = 39;
			IP[10] = 7;
			IP[11] = 47;
			IP[12] = 15;
			IP[13] = 55;
			IP[14] = 23;
			IP[15] = 63;
			IP[16] = 31;
			IP[17] = 38;
			IP[18] = 6;
			IP[19] = 46;
			IP[20] = 14;
			IP[21] = 54;
			IP[22] = 22;
			IP[23] = 62;
			IP[24] = 30;
			IP[25] = 37;
			IP[26] = 5;
			IP[27] = 45;
			IP[28] = 13;
			IP[29] = 53;
			IP[30] = 21;
			IP[31] = 61;
			IP[32] = 29;
			IP[33] = 36;
			IP[34] = 4;
			IP[35] = 44;
			IP[36] = 12;
			IP[37] = 52;
			IP[38] = 20;
			IP[39] = 60;
			IP[40] = 28;
			IP[41] = 35;
			IP[42] = 3;
			IP[43] = 43;
			IP[44] = 11;
			IP[45] = 51;
			IP[46] = 19;
			IP[47] = 59;
			IP[48] = 27;
			IP[49] = 34;
			IP[50] = 2;
			IP[51] = 42;
			IP[52] = 10;
			IP[53] = 50;
			IP[54] = 18;
			IP[55] = 58;
			IP[56] = 26;
			IP[57] = 33;
			IP[58] = 1;
			IP[59] = 41;
			IP[60] = 9;
			IP[61] = 49;
			IP[62] = 17;
			IP[63] = 57;
			IP[64] = 25;
              for(i=1; i<65; i++)
              z[i] = img[IP[i]];
              end
       endfunction

       function [48:1] exp(input [32:1] Ri);
        integer E[48:1];
        reg [48:1]z2;
        integer i;
              begin
                     E[1] = 32;
			E[2] = 1;
			E[3] = 2;
			E[4] = 3;
			E[5] = 4;
			E[6] = 5;
			E[7] = 4;
			E[8] = 5;
			E[9] = 6;
			E[10] = 7;
			E[11] = 8;
			E[12] = 9;
			E[13] = 8;
			E[14] = 9;
			E[15] = 10;
			E[16] = 11;
			E[17] = 12;
			E[18] = 13;
			E[19] = 12;
			E[20] = 13;
			E[21] = 14;
			E[22] = 15;
			E[23] = 16;
			E[24] = 17;
			E[25] = 16;
			E[26] = 17;
			E[27] = 18;
			E[28] = 19;
			E[29] = 20;
			E[30] = 21;
			E[31] = 20;
			E[32] = 21;
			E[33] = 22;
			E[34] = 23;
			E[35] = 24;
			E[36] = 25;
			E[37] = 24;
			E[38] = 25;
			E[39] = 26;
			E[40] = 27;
			E[41] = 28;
			E[42] = 29;
			E[43] = 28;
			E[44] = 29;
			E[45] = 30;
			E[46] = 31;
			E[47] = 32;
			E[48] = 1;
              for(i=1; i<49; i++)
              z2[i] = Ri[E[i]];
              end
       endfunction
       
       function [4:1] sub(input [6:1] sin,input n); // n is nth sub box
       integer s1[3:0][15:0] ;
       integer s2[3:0][15:0] ;
       integer s3[3:0][15:0] ;
       integer s4[3:0][15:0] ;
       integer s5[3:0][15:0] ;
       integer s6[3:0][15:0] ;
       integer s7[3:0][15:0] ;
       integer s8[3:0][15:0] ;
        reg [2:1] m;
        reg [4:1] l;
       begin
s1[0][0] = 14;s1[0][1] = 4;s1[0][2] = 13;s1[0][3] = 1;s1[0][4] = 2;s1[0][5] = 15;s1[0][6] = 11;s1[0][7] = 8;s1[0][8] = 3;s1[0][9] = 10;s1[0][10] = 6;s1[0][11] = 12;s1[0][12] = 5;s1[0][13] = 9;s1[0][14] = 0;s1[0][15] = 7;
s1[1][0] = 0;s1[1][1] = 15;s1[1][2] = 7;s1[1][3] = 4;s1[1][4] = 14;s1[1][5] = 2;s1[1][6] = 13;s1[1][7] = 1;s1[1][8] = 10;s1[1][9] = 6;s1[1][10] = 12;s1[1][11] = 11;s1[1][12] = 9;s1[1][13] = 5;s1[1][14] = 3;s1[1][15] = 8;
s1[2][0] = 4;s1[2][1] = 1;s1[2][2] = 14;s1[2][3] = 8;s1[2][4] = 13;s1[2][5] = 6;s1[2][6] = 2;s1[2][7] = 11;s1[2][8] = 15;s1[2][9] = 12;s1[2][10] = 9;s1[2][11] = 7;s1[2][12] = 3;s1[2][13] = 10;s1[2][14] = 5;s1[2][15] = 0;
s1[3][0] = 15;s1[3][1] = 12;s1[3][2] = 8;s1[3][3] = 2;s1[3][4] = 4;s1[3][5] = 9;s1[3][6] = 1;s1[3][7] = 7;s1[3][8] = 5;s1[3][9] = 11;s1[3][10] = 3;s1[3][11] = 14;s1[3][12] = 10;s1[3][13] = 0;s1[3][14] = 6;s1[3][15] = 13;
s2[0][0] = 15;s2[0][1] = 1;s2[0][2] = 8;s2[0][3] = 14;s2[0][4] = 6;s2[0][5] = 11;s2[0][6] = 3;s2[0][7] = 4;s2[0][8] = 9;s2[0][9] = 7;s2[0][10] = 2;s2[0][11] = 13;s2[0][12] = 12;s2[0][13] = 0;s2[0][14] = 5;s2[0][15] = 10;
s2[1][0] = 3;s2[1][1] = 13;s2[1][2] = 4;s2[1][3] = 7;s2[1][4] = 15;s2[1][5] = 2;s2[1][6] = 8;s2[1][7] = 14;s2[1][8] = 12;s2[1][9] = 0;s2[1][10] = 1;s2[1][11] = 10;s2[1][12] = 6;s2[1][13] = 9;s2[1][14] = 11;s2[1][15] = 5;
s2[2][0] = 0;s2[2][1] = 14;s2[2][2] = 7;s2[2][3] = 11;s2[2][4] = 10;s2[2][5] = 4;s2[2][6] = 13;s2[2][7] = 1;s2[2][8] = 5;s2[2][9] = 8;s2[2][10] = 12;s2[2][11] = 6;s2[2][12] = 9;s2[2][13] = 3;s2[2][14] = 2;s2[2][15] = 15;
s2[3][0] = 13;s2[3][1] = 8;s2[3][2] = 10;s2[3][3] = 1;s2[3][4] = 3;s2[3][5] = 15;s2[3][6] = 4;s2[3][7] = 2;s2[3][8] = 11;s2[3][9] = 6;s2[3][10] = 7;s2[3][11] = 12;s2[3][12] = 0;s2[3][13] = 5;s2[3][14] = 14;s2[3][15] = 9;
s3[0][0] = 10;s3[0][1] = 0;s3[0][2] = 9;s3[0][3] = 14;s3[0][4] = 6;s3[0][5] = 3;s3[0][6] = 15;s3[0][7] = 5;s3[0][8] = 1;s3[0][9] = 13;s3[0][10] = 12;s3[0][11] = 7;s3[0][12] = 11;s3[0][13] = 4;s3[0][14] = 2;s3[0][15] = 8;
s3[1][0] = 13;s3[1][1] = 7;s3[1][2] = 0;s3[1][3] = 9;s3[1][4] = 3;s3[1][5] = 4;s3[1][6] = 6;s3[1][7] = 10;s3[1][8] = 2;s3[1][9] = 8;s3[1][10] = 5;s3[1][11] = 14;s3[1][12] = 12;s3[1][13] = 11;s3[1][14] = 15;s3[1][15] = 1;
s3[2][0] = 13;s3[2][1] = 6;s3[2][2] = 4;s3[2][3] = 9;s3[2][4] = 8;s3[2][5] = 15;s3[2][6] = 3;s3[2][7] = 0;s3[2][8] = 11;s3[2][9] = 1;s3[2][10] = 2;s3[2][11] = 12;s3[2][12] = 5;s3[2][13] = 10;s3[2][14] = 14;s3[2][15] = 7;
s3[3][0] = 1;s3[3][1] = 10;s3[3][2] = 13;s3[3][3] = 0;s3[3][4] = 6;s3[3][5] = 9;s3[3][6] = 8;s3[3][7] = 7;s3[3][8] = 4;s3[3][9] = 15;s3[3][10] = 14;s3[3][11] = 3;s3[3][12] = 11;s3[3][13] = 5;s3[3][14] = 2;s3[3][15] = 12;
s4[0][0] = 7;s4[0][1] = 13;s4[0][2] = 14;s4[0][3] = 3;s4[0][4] = 0;s4[0][5] = 6;s4[0][6] = 9;s4[0][7] = 10;s4[0][8] = 1;s4[0][9] = 2;s4[0][10] = 8;s4[0][11] = 5;s4[0][12] = 11;s4[0][13] = 12;s4[0][14] = 4;s4[0][15] = 15;
s4[1][0] = 13;s4[1][1] = 8;s4[1][2] = 11;s4[1][3] = 5;s4[1][4] = 6;s4[1][5] = 15;s4[1][6] = 0;s4[1][7] = 3;s4[1][8] = 4;s4[1][9] = 7;s4[1][10] = 2;s4[1][11] = 12;s4[1][12] = 1;s4[1][13] = 10;s4[1][14] = 14;s4[1][15] = 9;
s4[2][0] = 10;s4[2][1] = 6;s4[2][2] = 9;s4[2][3] = 0;s4[2][4] = 12;s4[2][5] = 11;s4[2][6] = 7;s4[2][7] = 13;s4[2][8] = 15;s4[2][9] = 1;s4[2][10] = 3;s4[2][11] = 14;s4[2][12] = 5;s4[2][13] = 2;s4[2][14] = 8;s4[2][15] = 4;
s4[3][0] = 3;s4[3][1] = 15;s4[3][2] = 0;s4[3][3] = 6;s4[3][4] = 10;s4[3][5] = 1;s4[3][6] = 13;s4[3][7] = 8;s4[3][8] = 9;s4[3][9] = 4;s4[3][10] = 5;s4[3][11] = 11;s4[3][12] = 12;s4[3][13] = 7;s4[3][14] = 2;s4[3][15] = 14;
s5[0][0] = 2;s5[0][1] = 12;s5[0][2] = 4;s5[0][3] = 1;s5[0][4] = 7;s5[0][5] = 10;s5[0][6] = 11;s5[0][7] = 6;s5[0][8] = 8;s5[0][9] = 5;s5[0][10] = 3;s5[0][11] = 15;s5[0][12] = 13;s5[0][13] = 0;s5[0][14] = 14;s5[0][15] = 9;
s5[1][0] = 14;s5[1][1] = 11;s5[1][2] = 2;s5[1][3] = 12;s5[1][4] = 4;s5[1][5] = 7;s5[1][6] = 13;s5[1][7] = 1;s5[1][8] = 5;s5[1][9] = 0;s5[1][10] = 15;s5[1][11] = 10;s5[1][12] = 3;s5[1][13] = 9;s5[1][14] = 8;s5[1][15] = 6;
s5[2][0] = 4;s5[2][1] = 2;s5[2][2] = 1;s5[2][3] = 11;s5[2][4] = 10;s5[2][5] = 13;s5[2][6] = 7;s5[2][7] = 8;s5[2][8] = 15;s5[2][9] = 9;s5[2][10] = 12;s5[2][11] = 5;s5[2][12] = 6;s5[2][13] = 3;s5[2][14] = 0;s5[2][15] = 14;
s5[3][0] = 11;s5[3][1] = 8;s5[3][2] = 12;s5[3][3] = 7;s5[3][4] = 1;s5[3][5] = 14;s5[3][6] = 2;s5[3][7] = 13;s5[3][8] = 6;s5[3][9] = 15;s5[3][10] = 0;s5[3][11] = 9;s5[3][12] = 10;s5[3][13] = 4;s5[3][14] = 5;s5[3][15] = 3;
s6[0][0] = 12;s6[0][1] = 1;s6[0][2] = 10;s6[0][3] = 15;s6[0][4] = 9;s6[0][5] = 2;s6[0][6] = 6;s6[0][7] = 8;s6[0][8] = 0;s6[0][9] = 13;s6[0][10] = 3;s6[0][11] = 4;s6[0][12] = 14;s6[0][13] = 7;s6[0][14] = 5;s6[0][15] = 11;
s6[1][0] = 10;s6[1][1] = 15;s6[1][2] = 4;s6[1][3] = 2;s6[1][4] = 7;s6[1][5] = 12;s6[1][6] = 9;s6[1][7] = 5;s6[1][8] = 6;s6[1][9] = 1;s6[1][10] = 13;s6[1][11] = 14;s6[1][12] = 0;s6[1][13] = 11;s6[1][14] = 3;s6[1][15] = 8;
s6[2][0] = 9;s6[2][1] = 14;s6[2][2] = 15;s6[2][3] = 5;s6[2][4] = 2;s6[2][5] = 8;s6[2][6] = 12;s6[2][7] = 3;s6[2][8] = 7;s6[2][9] = 0;s6[2][10] = 4;s6[2][11] = 10;s6[2][12] = 1;s6[2][13] = 13;s6[2][14] = 11;s6[2][15] = 6;
s6[3][0] = 4;s6[3][1] = 3;s6[3][2] = 2;s6[3][3] = 12;s6[3][4] = 9;s6[3][5] = 5;s6[3][6] = 15;s6[3][7] = 10;s6[3][8] = 11;s6[3][9] = 14;s6[3][10] = 1;s6[3][11] = 7;s6[3][12] = 6;s6[3][13] = 0;s6[3][14] = 8;s6[3][15] = 13;
s7[0][0] = 4;s7[0][1] = 11;s7[0][2] = 2;s7[0][3] = 14;s7[0][4] = 15;s7[0][5] = 0;s7[0][6] = 8;s7[0][7] = 13;s7[0][8] = 3;s7[0][9] = 12;s7[0][10] = 9;s7[0][11] = 7;s7[0][12] = 5;s7[0][13] = 10;s7[0][14] = 6;s7[0][15] = 1;
s7[1][0] = 13;s7[1][1] = 0;s7[1][2] = 11;s7[1][3] = 7;s7[1][4] = 4;s7[1][5] = 9;s7[1][6] = 1;s7[1][7] = 10;s7[1][8] = 14;s7[1][9] = 3;s7[1][10] = 5;s7[1][11] = 12;s7[1][12] = 2;s7[1][13] = 15;s7[1][14] = 8;s7[1][15] = 6;
s7[2][0] = 1;s7[2][1] = 4;s7[2][2] = 11;s7[2][3] = 13;s7[2][4] = 12;s7[2][5] = 3;s7[2][6] = 7;s7[2][7] = 14;s7[2][8] = 10;s7[2][9] = 15;s7[2][10] = 6;s7[2][11] = 8;s7[2][12] = 0;s7[2][13] = 5;s7[2][14] = 9;s7[2][15] = 2;
s7[3][0] = 6;s7[3][1] = 11;s7[3][2] = 13;s7[3][3] = 8;s7[3][4] = 1;s7[3][5] = 4;s7[3][6] = 10;s7[3][7] = 7;s7[3][8] = 9;s7[3][9] = 5;s7[3][10] = 0;s7[3][11] = 15;s7[3][12] = 14;s7[3][13] = 2;s7[3][14] = 3;s7[3][15] = 12;
s8[0][0] = 13;s8[0][1] = 2;s8[0][2] = 8;s8[0][3] = 4;s8[0][4] = 6;s8[0][5] = 15;s8[0][6] = 11;s8[0][7] = 1;s8[0][8] = 10;s8[0][9] = 9;s8[0][10] = 3;s8[0][11] = 14;s8[0][12] = 5;s8[0][13] = 0;s8[0][14] = 12;s8[0][15] = 7;
s8[1][0] = 1;s8[1][1] = 15;s8[1][2] = 13;s8[1][3] = 8;s8[1][4] = 10;s8[1][5] = 3;s8[1][6] = 7;s8[1][7] = 4;s8[1][8] = 12;s8[1][9] = 5;s8[1][10] = 6;s8[1][11] = 11;s8[1][12] = 0;s8[1][13] = 14;s8[1][14] = 9;s8[1][15] = 2;
s8[2][0] = 7;s8[2][1] = 11;s8[2][2] = 4;s8[2][3] = 1;s8[2][4] = 9;s8[2][5] = 12;s8[2][6] = 14;s8[2][7] = 2;s8[2][8] = 0;s8[2][9] = 6;s8[2][10] = 10;s8[2][11] = 13;s8[2][12] = 15;s8[2][13] = 3;s8[2][14] = 5;s8[2][15] = 8;
s8[3][0] = 2;s8[3][1] = 1;s8[3][2] = 14;s8[3][3] = 7;s8[3][4] = 4;s8[3][5] = 10;s8[3][6] = 8;s8[3][7] = 13;s8[3][8] = 15;s8[3][9] = 12;s8[3][10] = 9;s8[3][11] = 0;s8[3][12] = 3;s8[3][13] = 5;s8[3][14] = 6;s8[3][15] = 11;
       m[2:1] = {sin[6], sin[1]};
       l[4:1] = sin[5:2];
                  
        case(n)
        4'b0001:sub = s1[m][l];
        4'b0010:sub = s1[m][l];
        4'b0011:sub = s1[m][l];
        4'b0010:sub = s1[m][l];
        4'b0010:sub = s1[m][l];
        4'b0010:sub = s1[m][l];
        endcase
                    end
       endfunction
        
       
       function [32:1] perm_P(input [32:1] s_res);
     integer i;
     integer P[32:1];
     reg [32:1] temp_P;
     begin
		       P[1] = 16;
			P[2] = 7;
			P[3] = 20;
			P[4] = 21;
			P[5] = 29;
			P[6] = 12;
			P[7] = 28;
			P[8] = 17;
			P[9] = 1;
			P[10] = 15;
			P[11] = 23;
			P[12] = 26;
			P[13] = 5;
			P[14] = 18;
			P[15] = 31;
			P[16] = 10;
			P[17] = 2;
			P[18] = 8;
			P[19] = 24;
			P[20] = 14;
			P[21] = 32;
			P[22] = 27;
			P[23] = 3;
			P[24] = 9;
			P[25] = 19;
			P[26] = 13;
			P[27] = 30;
			P[28] = 6;
			P[29] = 22;
			P[30] = 11;
			P[31] = 4;
			P[32] = 25;

      for(i=1; i<=32; i=i+1)
      temp_P[32-i+1] = s_res[32-P[i]+1];
      perm_P = temp_P;
    end
  endfunction
       

function [64:1] IPinverse(input [64:1] message);
	  integer IPin[64:1];
     reg [64:1] temp_msg;
     integer i;
 	  begin
			IPin[1] = 40;
			IPin[2] = 8;
			IPin[3] = 48;
			IPin[4] = 16;
			IPin[5] = 56;
			IPin[6] = 24;
			IPin[7] = 64;
			IPin[8] = 32;
			IPin[9] = 39;
			IPin[10] = 7;
			IPin[11] = 47;
			IPin[12] = 15;
			IPin[13] = 55;
			IPin[14] = 23;
			IPin[15] = 63;
			IPin[16] = 31;
			IPin[17] = 38;
			IPin[18] = 6;
			IPin[19] = 46;
			IPin[20] = 14;
			IPin[21] = 54;
			IPin[22] = 22;
			IPin[23] = 62;
			IPin[24] = 30;
			IPin[25] = 37;
			IPin[26] = 5;
			IPin[27] = 45;
			IPin[28] = 13;
			IPin[29] = 53;
			IPin[30] = 21;
			IPin[31] = 61;
			IPin[32] = 29;
			IPin[33] = 36;
			IPin[34] = 4;
			IPin[35] = 44;
			IPin[36] = 12;
			IPin[37] = 52;
			IPin[38] = 20;
			IPin[39] = 60;
			IPin[40] = 28;
			IPin[41] = 35;
			IPin[42] = 3;
			IPin[43] = 43;
			IPin[44] = 11;
			IPin[45] = 51;
			IPin[46] = 19;
			IPin[47] = 59;
			IPin[48] = 27;
			IPin[49] = 34;
			IPin[50] = 2;
			IPin[51] = 42;
			IPin[52] = 10;
			IPin[53] = 50;
			IPin[54] = 18;
			IPin[55] = 58;
			IPin[56] = 26;
			IPin[57] = 33;
			IPin[58] = 1;
			IPin[59] = 41;
			IPin[60] = 9;
			IPin[61] = 49;
			IPin[62] = 17;
			IPin[63] = 57;
			IPin[64] = 25;

			for(i=1; i<=64; i=i+1)
            temp_msg[i] = message[IPin[i]];
           IPinverse = temp_msg;
 	  end
  endfunction
       
    function [32:1] f(input [32:1] R, input [48:1] K);
    reg [48:1] temp;
    reg [32:1] temp_after_s_box;
    reg [5:0] B[8:1];
    begin
      temp = K ^ exp(R);
      B[1] = temp[48:43];
      B[2] = temp[42:37];
      B[3] = temp[36:31];
      B[4] = temp[30:25];
      B[5] = temp[24:19];
      B[6] = temp[18:13];
      B[7] = temp[12:7];
      B[8] = temp[6:1];
      
      temp_after_s_box = {sub(B[1], 5'd1), sub(B[2], 5'd2), sub(B[3], 5'd3), sub(B[4], 5'd4),
                          sub(B[5], 5'd5), sub(B[6], 5'd6), sub(B[7], 5'd7), sub(B[8], 5'd8)};

      f = perm_P(temp_after_s_box);
    end
  endfunction    

  reg [64:1] new_msg;
  reg [32:1] L[16:0], R[16:0];
  wire [48:1] k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15, k16;
  reg [48:1] K[16:1];
  integer i;
  ProcessKey pk(k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15, k16, key);

  always @(*)
  begin
    new_msg = IPerm(img);
    {L[0], R[0]} = new_msg;

    K[1] = k1; K[2] = k2; K[3] = k3; K[4] = k4; K[5] = k5; K[6] = k6; K[7] = k7; K[8] = k8; K[9] = k9; K[10] = k10; K[11] = k11; K[12] = k12; K[13] = k13; K[14] = k14; K[15] = k15; K[16] = k16; 

    for(i=1; i<=16; i=i+1)
    begin
      L[i]=R[i-1];
      R[i]=L[i-1] ^ f(R[i-1], K[i]);
    end
    enigma[64:1] = IPinverse({R[16], L[16]});
  end  
endmodule
